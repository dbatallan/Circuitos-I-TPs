** Profile: "SCHEMATIC1-ACanalysis"  [ C:\Users\Lionheart\Documents\GitHub\Circuitos-I-TPs\TL2\Simulaciones\Monoetapa\JFETN\PSPICE\JFETN-PSpiceFiles\SCHEMATIC1\ACanalysis.sim ] 

** Creating circuit file "ACanalysis.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 30 1 100Meg
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
